library verilog;
use verilog.vl_types.all;
entity ekf is
    generic(
        SIGN            : integer := 1;
        INT_CASE1       : integer := 0;
        FR_CASE1        : integer := 23;
        INT_CASE2       : integer := 2;
        FR_CASE2        : integer := 21;
        INT_CASE3       : integer := 7;
        FR_CASE3        : integer := 16;
        D_WIDTH         : integer := 24;
        STATE_CNT       : integer := 3;
        IDLE            : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi0);
        LATENCY_1       : vl_logic_vector(0 to 2) := (Hi0, Hi0, Hi1);
        LATENCY_2       : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi0);
        LATENCY_3       : vl_logic_vector(0 to 2) := (Hi0, Hi1, Hi1);
        LATENCY_4       : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi0);
        LATENCY_5       : vl_logic_vector(0 to 2) := (Hi1, Hi0, Hi1);
        DONE            : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi0);
        SOC_DONE        : vl_logic_vector(0 to 2) := (Hi1, Hi1, Hi1);
        RI              : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1);
        RD              : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        CD              : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1);
        CB              : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1);
        Q_1             : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        Q_4             : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        R               : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        b_1_1000        : vl_logic_vector(0 to 23) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        b_2_1000        : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        a_4_1000        : vl_logic_vector(0 to 23) := (Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0);
        a_4_1000_2      : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        b_1_100         : vl_logic_vector(0 to 23) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0);
        b_2_100         : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1);
        a_4_100         : vl_logic_vector(0 to 23) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0);
        a_4_100_2       : vl_logic_vector(0 to 23) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        theta4_1        : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0);
        theta4_2        : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0);
        theta4_3        : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1);
        theta5_1        : vl_logic_vector(0 to 23) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        theta5_2        : vl_logic_vector(0 to 23) := (Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        theta5_3        : vl_logic_vector(0 to 23) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        dt_cd_ri_1000   : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi1, Hi1);
        dt_cd_ri_100    : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        first_p1        : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        first_p2        : vl_notype;
        first_p3        : vl_notype;
        first_p4        : vl_logic_vector(0 to 23) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0)
    );
    port(
        clk             : in     vl_logic;
        n_rst           : in     vl_logic;
        start           : in     vl_logic;
        ekf_vrc         : out    vl_logic_vector;
        ekf_soc         : out    vl_logic_vector;
        ekf_done        : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of SIGN : constant is 1;
    attribute mti_svvh_generic_type of INT_CASE1 : constant is 1;
    attribute mti_svvh_generic_type of FR_CASE1 : constant is 1;
    attribute mti_svvh_generic_type of INT_CASE2 : constant is 1;
    attribute mti_svvh_generic_type of FR_CASE2 : constant is 1;
    attribute mti_svvh_generic_type of INT_CASE3 : constant is 1;
    attribute mti_svvh_generic_type of FR_CASE3 : constant is 1;
    attribute mti_svvh_generic_type of D_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of STATE_CNT : constant is 1;
    attribute mti_svvh_generic_type of IDLE : constant is 1;
    attribute mti_svvh_generic_type of LATENCY_1 : constant is 1;
    attribute mti_svvh_generic_type of LATENCY_2 : constant is 1;
    attribute mti_svvh_generic_type of LATENCY_3 : constant is 1;
    attribute mti_svvh_generic_type of LATENCY_4 : constant is 1;
    attribute mti_svvh_generic_type of LATENCY_5 : constant is 1;
    attribute mti_svvh_generic_type of DONE : constant is 1;
    attribute mti_svvh_generic_type of SOC_DONE : constant is 1;
    attribute mti_svvh_generic_type of RI : constant is 1;
    attribute mti_svvh_generic_type of RD : constant is 1;
    attribute mti_svvh_generic_type of CD : constant is 1;
    attribute mti_svvh_generic_type of CB : constant is 1;
    attribute mti_svvh_generic_type of Q_1 : constant is 1;
    attribute mti_svvh_generic_type of Q_4 : constant is 1;
    attribute mti_svvh_generic_type of R : constant is 1;
    attribute mti_svvh_generic_type of b_1_1000 : constant is 1;
    attribute mti_svvh_generic_type of b_2_1000 : constant is 1;
    attribute mti_svvh_generic_type of a_4_1000 : constant is 1;
    attribute mti_svvh_generic_type of a_4_1000_2 : constant is 1;
    attribute mti_svvh_generic_type of b_1_100 : constant is 1;
    attribute mti_svvh_generic_type of b_2_100 : constant is 1;
    attribute mti_svvh_generic_type of a_4_100 : constant is 1;
    attribute mti_svvh_generic_type of a_4_100_2 : constant is 1;
    attribute mti_svvh_generic_type of theta4_1 : constant is 1;
    attribute mti_svvh_generic_type of theta4_2 : constant is 1;
    attribute mti_svvh_generic_type of theta4_3 : constant is 1;
    attribute mti_svvh_generic_type of theta5_1 : constant is 1;
    attribute mti_svvh_generic_type of theta5_2 : constant is 1;
    attribute mti_svvh_generic_type of theta5_3 : constant is 1;
    attribute mti_svvh_generic_type of dt_cd_ri_1000 : constant is 1;
    attribute mti_svvh_generic_type of dt_cd_ri_100 : constant is 1;
    attribute mti_svvh_generic_type of first_p1 : constant is 1;
    attribute mti_svvh_generic_type of first_p2 : constant is 3;
    attribute mti_svvh_generic_type of first_p3 : constant is 3;
    attribute mti_svvh_generic_type of first_p4 : constant is 1;
end ekf;
